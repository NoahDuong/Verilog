----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:36:49 09/23/2024 
-- Design Name: 
-- Module Name:    UPDOWNCOUNTER - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity UPDOWNCOUNTER is
    Port ( Clk : in  STD_LOGIC;
           RST : in  STD_LOGIC;
           OUT : out  STD_LOGIC_VECTOR (3 downto 0));
end UPDOWNCOUNTER;

architecture Behavioral of UPDOWNCOUNTER is

begin


end Behavioral;

